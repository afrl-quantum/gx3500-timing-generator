// megafunction wizard: %ALTIOBUF%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altiobuf_out 

// ============================================================
// File Name: Driver128b.v
// Megafunction Name(s):
// 			altiobuf_out
//
// Simulation Library Files(s):
// 			cycloneiii
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.0 Build 162 10/23/2013 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module Driver128b (
	datain,
	dataout)/* synthesis synthesis_clearbox = 1 */;

	input	[127:0]  datain;
	output	[127:0]  dataout;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
// Retrieval info: CONSTANT: left_shift_series_termination_control STRING "FALSE"
// Retrieval info: CONSTANT: number_of_channels NUMERIC "128"
// Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
// Retrieval info: CONSTANT: pseudo_differential_mode STRING "FALSE"
// Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
// Retrieval info: CONSTANT: use_oe STRING "FALSE"
// Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
// Retrieval info: USED_PORT: datain 0 0 128 0 INPUT NODEFVAL "datain[127..0]"
// Retrieval info: USED_PORT: dataout 0 0 128 0 OUTPUT NODEFVAL "dataout[127..0]"
// Retrieval info: CONNECT: @datain 0 0 128 0 datain 0 0 128 0
// Retrieval info: CONNECT: dataout 0 0 128 0 @dataout 0 0 128 0
// Retrieval info: GEN_FILE: TYPE_NORMAL Driver128b.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Driver128b.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Driver128b.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Driver128b.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Driver128b_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Driver128b_bb.v TRUE
// Retrieval info: LIB_FILE: cycloneiii
