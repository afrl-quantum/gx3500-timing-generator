// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Thu Aug 13 11:50:28 2015

// synthesis message_off 10175

`timescale 1ns/1ns

module System_State (
    reset,clock,Do_Arm,Do_Stop,Do_Trigger,PCI_Enabled,Buffer_Empty,Do_Repeat,Do_Pause,Do_Resume,Is_Finished,
    PCI_Allowed,Internal_State[2:0],Load_Instructions,Run_Timer,Reset_Timer,Output_Sequence);

    input reset;
    input clock;
    input Do_Arm;
    input Do_Stop;
    input Do_Trigger;
    input PCI_Enabled;
    input Buffer_Empty;
    input Do_Repeat;
    input Do_Pause;
    input Do_Resume;
    input Is_Finished;
    tri0 reset;
    tri0 Do_Arm;
    tri0 Do_Stop;
    tri0 Do_Trigger;
    tri0 PCI_Enabled;
    tri0 Buffer_Empty;
    tri0 Do_Repeat;
    tri0 Do_Pause;
    tri0 Do_Resume;
    tri0 Is_Finished;
    output PCI_Allowed;
    output [2:0] Internal_State;
    output Load_Instructions;
    output Run_Timer;
    output Reset_Timer;
    output Output_Sequence;
    reg PCI_Allowed;
    reg [2:0] Internal_State;
    reg Load_Instructions;
    reg Run_Timer;
    reg Reset_Timer;
    reg Output_Sequence;
    reg [6:0] fstate;
    reg [6:0] reg_fstate;
    parameter STOPPING=0,ARMING1=1,READY=2,SETUP=3,ARMING2=4,RUN=5,PAUSED=6;

    always @(posedge clock or negedge reset)
    begin
        if (~reset) begin
            fstate <= STOPPING;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or Do_Arm or Do_Stop or Do_Trigger or PCI_Enabled or Buffer_Empty or Do_Repeat or Do_Pause or Do_Resume or Is_Finished)
    begin
        PCI_Allowed <= 1'b0;
        Internal_State <= 3'b000;
        Load_Instructions <= 1'b0;
        Run_Timer <= 1'b0;
        Reset_Timer <= 1'b0;
        Output_Sequence <= 1'b0;
        case (fstate)
            STOPPING: begin
                if (PCI_Enabled)
                    reg_fstate <= SETUP;
                else if (~(PCI_Enabled))
                    reg_fstate <= STOPPING;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= STOPPING;

                Output_Sequence <= 1'b0;

                Internal_State <= 3'b101;

                PCI_Allowed <= 1'b1;

                Reset_Timer <= 1'b0;

                Run_Timer <= 1'b0;

                Load_Instructions <= 1'b0;
            end
            ARMING1: begin
                if (~(PCI_Enabled))
                    reg_fstate <= ARMING2;
                else if (PCI_Enabled)
                    reg_fstate <= ARMING1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= ARMING1;

                Output_Sequence <= 1'b0;

                Internal_State <= 3'b100;

                PCI_Allowed <= 1'b0;

                Reset_Timer <= 1'b1;

                Run_Timer <= 1'b0;

                Load_Instructions <= 1'b0;
            end
            READY: begin
                if ((Do_Trigger & ~(Do_Stop)))
                    reg_fstate <= RUN;
                else if (Do_Stop)
                    reg_fstate <= STOPPING;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= READY;

                Output_Sequence <= 1'b0;

                Internal_State <= 3'b001;

                PCI_Allowed <= 1'b0;

                Reset_Timer <= 1'b0;

                Run_Timer <= 1'b0;

                Load_Instructions <= 1'b1;
            end
            SETUP: begin
                if (Do_Arm)
                    reg_fstate <= ARMING1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= SETUP;

                Output_Sequence <= 1'b0;

                Internal_State <= 3'b000;

                PCI_Allowed <= 1'b1;

                Reset_Timer <= 1'b0;

                Run_Timer <= 1'b0;

                Load_Instructions <= 1'b0;
            end
            ARMING2: begin
                if (~(Buffer_Empty))
                    reg_fstate <= READY;
                else if (Buffer_Empty)
                    reg_fstate <= ARMING2;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= ARMING2;

                Output_Sequence <= 1'b0;

                Internal_State <= 3'b100;

                PCI_Allowed <= 1'b0;

                Reset_Timer <= 1'b0;

                Run_Timer <= 1'b0;

                Load_Instructions <= 1'b1;
            end
            RUN: begin
                if ((Do_Repeat & ~(((Do_Stop | Is_Finished) | Do_Pause))))
                    reg_fstate <= ARMING1;
                else if ((Do_Pause & ~((Do_Stop | Is_Finished))))
                    reg_fstate <= PAUSED;
                else if ((Do_Stop | Is_Finished))
                    reg_fstate <= STOPPING;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= RUN;

                Output_Sequence <= 1'b1;

                Internal_State <= 3'b010;

                PCI_Allowed <= 1'b0;

                Reset_Timer <= 1'b0;

                Run_Timer <= 1'b1;

                Load_Instructions <= 1'b1;
            end
            PAUSED: begin
                if ((Do_Resume & ~(Do_Stop)))
                    reg_fstate <= RUN;
                else if (Do_Stop)
                    reg_fstate <= STOPPING;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= PAUSED;

                Output_Sequence <= 1'b1;

                Internal_State <= 3'b011;

                PCI_Allowed <= 1'b0;

                Reset_Timer <= 1'b0;

                Run_Timer <= 1'b0;

                Load_Instructions <= 1'b1;
            end
            default: begin
                PCI_Allowed <= 1'bx;
                Internal_State <= 3'bxxx;
                Load_Instructions <= 1'bx;
                Run_Timer <= 1'bx;
                Reset_Timer <= 1'bx;
                Output_Sequence <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // System_State
