// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Wed Aug 12 11:33:33 2015

// synthesis message_off 10175

`timescale 1ns/1ns

module RAM_Clock_Switch (
    reset,clock,PCI_Allowed,
    UsePCI,PCI_Enabled,RAM_Enabled,UsePCIClock);

    input reset;
    input clock;
    input PCI_Allowed;
    tri0 reset;
    tri0 PCI_Allowed;
    output UsePCI;
    output PCI_Enabled;
    output RAM_Enabled;
    output UsePCIClock;
    reg UsePCI;
    reg PCI_Enabled;
    reg RAM_Enabled;
    reg UsePCIClock;
    reg [16:0] fstate;
    reg [16:0] reg_fstate;
    parameter NoPCI_RAM_Disabled_L=0,PCI_RAM_Disabled_L=1,Steady_State_NoPCI=2,Start=3,Steady_State_PCI=4,PCI_RAM_Disabled_R=5,NoPCI_RAM_Disabled_R=6,RWait1=7,RWait2=8,RWait3=9,RWait4=10,LWait1=11,LWait2=12,LWait3=13,LWait4=14,NoPCI_Clock=15,PCI_Clock=16;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or PCI_Allowed)
    begin
        if (~reset) begin
            reg_fstate <= Start;
            UsePCI <= 1'b0;
            PCI_Enabled <= 1'b0;
            RAM_Enabled <= 1'b0;
            UsePCIClock <= 1'b0;
        end
        else begin
            UsePCI <= 1'b0;
            PCI_Enabled <= 1'b0;
            RAM_Enabled <= 1'b0;
            UsePCIClock <= 1'b0;
            case (fstate)
                NoPCI_RAM_Disabled_L: begin
                    reg_fstate <= LWait1;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b0;
                end
                PCI_RAM_Disabled_L: begin
                    reg_fstate <= PCI_Clock;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b0;
                end
                Steady_State_NoPCI: begin
                    if (PCI_Allowed)
                        reg_fstate <= NoPCI_RAM_Disabled_L;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Steady_State_NoPCI;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b1;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b0;
                end
                Start: begin
                    if (PCI_Allowed)
                        reg_fstate <= NoPCI_RAM_Disabled_L;
                    else if (~(PCI_Allowed))
                        reg_fstate <= PCI_RAM_Disabled_R;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Start;

                    PCI_Enabled <= PCI_Allowed;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= PCI_Allowed;

                    UsePCIClock <= PCI_Allowed;
                end
                Steady_State_PCI: begin
                    if (~(PCI_Allowed))
                        reg_fstate <= PCI_RAM_Disabled_R;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Steady_State_PCI;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b1;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b1;
                end
                PCI_RAM_Disabled_R: begin
                    reg_fstate <= RWait1;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b1;
                end
                NoPCI_RAM_Disabled_R: begin
                    reg_fstate <= NoPCI_Clock;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b1;
                end
                RWait1: begin
                    reg_fstate <= RWait2;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b1;
                end
                RWait2: begin
                    reg_fstate <= NoPCI_RAM_Disabled_R;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b1;
                end
                RWait3: begin
                    reg_fstate <= RWait4;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b0;
                end
                RWait4: begin
                    reg_fstate <= Steady_State_NoPCI;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b0;
                end
                LWait1: begin
                    reg_fstate <= LWait2;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b0;
                end
                LWait2: begin
                    reg_fstate <= PCI_RAM_Disabled_L;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b0;
                end
                LWait3: begin
                    reg_fstate <= LWait4;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b1;
                end
                LWait4: begin
                    reg_fstate <= Steady_State_PCI;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b1;
                end
                NoPCI_Clock: begin
                    reg_fstate <= RWait3;

                    PCI_Enabled <= 1'b1;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b0;

                    UsePCIClock <= 1'b0;
                end
                PCI_Clock: begin
                    reg_fstate <= LWait3;

                    PCI_Enabled <= 1'b0;

                    RAM_Enabled <= 1'b0;

                    UsePCI <= 1'b1;

                    UsePCIClock <= 1'b1;
                end
                default: begin
                    UsePCI <= 1'bx;
                    PCI_Enabled <= 1'bx;
                    RAM_Enabled <= 1'bx;
                    UsePCIClock <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // RAM_Clock_Switch
